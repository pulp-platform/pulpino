
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h81868106,
    32'h82868206,
    32'h83868306,
    32'h84868406,
    32'h85868506,
    32'h86868606,
    32'h87868706,
    32'h88868806,
    32'h89868906,
    32'h8A868A06,
    32'h8B868B06,
    32'h8C868C06,
    32'h8D868D06,
    32'h8E868E06,
    32'h8F868F06,
    32'h00100117,
    32'hF3010113,
    32'h00000D17,
    32'h5B8D0D13,
    32'h00000D97,
    32'h5B0D8D93,
    32'h01BD5763,
    32'h000D2023,
    32'hDDE30D11,
    32'h0513FFAD,
    32'h05930000,
    32'h00EF0000,
    32'h00000740,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h11010000,
    32'h46014681,
    32'h051345A1,
    32'hCE0609F0,
    32'h348000EF,
    32'h04000513,
    32'h378000EF,
    32'h45014581,
    32'h360000EF,
    32'h45014581,
    32'h388000EF,
    32'h05930028,
    32'h00EF0400,
    32'h47A23B20,
    32'h21900713,
    32'h0187D513,
    32'h157D87A1,
    32'h1007D7B3,
    32'h00A03533,
    32'h00E78863,
    32'h07616709,
    32'h37B38F99,
    32'h953E00F0,
    32'h610540F2,
    32'h715D8082,
    32'hC6864505,
    32'hC2A6C4A2,
    32'hDE4EC0CA,
    32'hDA56DC52,
    32'hD65ED85A,
    32'hD266D462,
    32'h00EFD06A,
    32'h45852660,
    32'h00EF4501,
    32'h67853AA0,
    32'hBB878793,
    32'h0037C0FB,
    32'h00010001,
    32'h27B74711,
    32'hC3D81A10,
    32'hF63FF0EF,
    32'h8537C911,
    32'h05930000,
    32'h05130240,
    32'h00EF5E85,
    32'hA0013BA0,
    32'h00008537,
    32'h051345C5,
    32'h00EF6105,
    32'h46813AA0,
    32'h45A14601,
    32'h00EF4519,
    32'h450128A0,
    32'h2BC000EF,
    32'h458164C1,
    32'h00EF4505,
    32'h14FD2D20,
    32'h00EF4405,
    32'h8D652EE0,
    32'hFE851DE3,
    32'h80000637,
    32'h02000693,
    32'h34860613,
    32'h051345A1,
    32'h00EF0710,
    32'h45012560,
    32'h288000EF,
    32'h458164C1,
    32'h00EF8522,
    32'h14FD29E0,
    32'h2BC000EF,
    32'h1DE38D65,
    32'h4581FE85,
    32'h00EF4521,
    32'h069325A0,
    32'h46010200,
    32'h051345A1,
    32'h00EF0EB0,
    32'h05132220,
    32'h00EF1000,
    32'h45812520,
    32'h00EF4509,
    32'h059326A0,
    32'h850A1000,
    32'h294000EF,
    32'h85374CB2,
    32'h45D50000,
    32'h62450513,
    32'h4C124402,
    32'h4AD249C2,
    32'h00EF4B72,
    32'h45813020,
    32'h00EF4521,
    32'h5F6320E0,
    32'h84A20790,
    32'h49016421,
    32'h409C0C33,
    32'h00008BB7,
    32'h68040413,
    32'h00008A37,
    32'h96136D05,
    32'h06930084,
    32'h45A10200,
    32'h0EB00513,
    32'h1B8000EF,
    32'h00EF6521,
    32'h45811EA0,
    32'h00EF4509,
    32'h05332020,
    32'h65A1009C,
    32'h22C000EF,
    32'h85134599,
    32'h00EF63CB,
    32'h55132AA0,
    32'h45850049,
    32'h00EF9522,
    32'h751329E0,
    32'h458500F9,
    32'h00EF9522,
    32'h09052920,
    32'h05134599,
    32'h00EF644A,
    32'h94EA2860,
    32'h2AC000EF,
    32'hFB2C91E3,
    32'h147D6441,
    32'h00EF4485,
    32'h8D611DA0,
    32'hFE951DE3,
    32'h00008537,
    32'h051345B5,
    32'h00EF64C5,
    32'h00EF25E0,
    32'h45812860,
    32'h00EF4521,
    32'h5F631660,
    32'h64210760,
    32'h490184CE,
    32'h413A89B3,
    32'h00008BB7,
    32'h68040413,
    32'h00008A37,
    32'h96136A85,
    32'h06930084,
    32'h45A10200,
    32'h0EB00513,
    32'h110000EF,
    32'h00EF6521,
    32'h45811420,
    32'h00EF4509,
    32'h853315A0,
    32'h65A10099,
    32'h184000EF,
    32'h85134599,
    32'h00EF63CB,
    32'h55132020,
    32'h45850049,
    32'h00EF9522,
    32'h75131F60,
    32'h458500F9,
    32'h00EF9522,
    32'h09051EA0,
    32'h05134599,
    32'h00EF644A,
    32'h94D61DE0,
    32'h204000EF,
    32'hFB2B11E3,
    32'h00008537,
    32'h02200593,
    32'h65C50513,
    32'h1C4000EF,
    32'h1EC000EF,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000793,
    32'h00078067,
    32'h00010001,
    32'h40B60001,
    32'h44264501,
    32'h49064496,
    32'h5A6259F2,
    32'h5B425AD2,
    32'h5C225BB2,
    32'h5D025C92,
    32'h80826161,
    32'hC4221141,
    32'h842A4581,
    32'hC606453D,
    32'h00EFC226,
    32'h45811B60,
    32'h00EF4539,
    32'h45811AE0,
    32'h00EF4535,
    32'h45811A60,
    32'h00EF4531,
    32'h5F6319E0,
    32'h44850280,
    32'h45414581,
    32'h190000EF,
    32'h02940863,
    32'h452D4581,
    32'h184000EF,
    32'h01634789,
    32'h458102F4,
    32'h00EF4501,
    32'h478D1760,
    32'h00F40A63,
    32'h40B28526,
    32'h44924422,
    32'h01414581,
    32'h1600006F,
    32'h442240B2,
    32'h01414492,
    32'h00008082,
    32'h07136711,
    32'h06A2F007,
    32'h02000793,
    32'h8EF98F8D,
    32'h03F5F593,
    32'h1A102737,
    32'h00F51533,
    32'hC7088DD5,
    32'hCB0CC750,
    32'h00008082,
    32'h553305C2,
    32'h8DC91005,
    32'h1A1027B7,
    32'h8082CBCC,
    32'h1A102737,
    32'h11414B1C,
    32'hC63E0542,
    32'hD7B347B2,
    32'h8D5D1007,
    32'h47B2C62A,
    32'hCB1C0141,
    32'h00008082,
    32'h05A14785,
    32'h00B795B3,
    32'h00A79533,
    32'h87936785,
    32'h8DFDF007,
    32'h0FF57513,
    32'h27B78D4D,
    32'hC3881A10,
    32'h00008082,
    32'h1A1027B7,
    32'h1141439C,
    32'h4532C63E,
    32'h80820141,
    32'h4055D793,
    32'hF7931141,
    32'h89FD7FF7,
    32'hC581C43E,
    32'h078547A2,
    32'hC602C43E,
    32'h47A246B2,
    32'h1A102737,
    32'hD36385BA,
    32'h431C02F6,
    32'hF79387C1,
    32'hDFE50FF7,
    32'h519046B2,
    32'h068A47B2,
    32'h1AC56023,
    32'hC63E0785,
    32'h47A246B2,
    32'hFEF6C1E3,
    32'h80820141,
    32'h1A1076B7,
    32'h07B742D8,
    32'hD6131A10,
    32'h67130085,
    32'hC2D80027,
    32'h08300713,
    32'hF593C7D8,
    32'h07130FF5,
    32'hC3D00A70,
    32'hC798C38C,
    32'hC7D8470D,
    32'h771343D8,
    32'h67130F07,
    32'hC3D80027,
    32'h00008082,
    32'h1A100737,
    32'h0693C185,
    32'h4B5C0400,
    32'h0207F793,
    32'h460BDFED,
    32'h07B70015,
    32'h15FD1A10,
    32'h16FDC390,
    32'hF1F5E299,
    32'hF1F58082,
    32'h00008082,
    32'h1A100737,
    32'hF7934B5C,
    32'hDFED0407,
    32'h00008082,
    32'h1A1076B7,
    32'h1141429C,
    32'h00A595B3,
    32'h4732C63E,
    32'h97B34785,
    32'hC79300A7,
    32'h8FF9FFF7,
    32'h47B2C63E,
    32'h00F5E533,
    32'h47B2C62A,
    32'hC29C0141,
    32'h00008082,
    32'h4F525245,
    32'h53203A52,
    32'h736E6170,
    32'h206E6F69,
    32'h20495053,
    32'h73616C66,
    32'h6F6E2068,
    32'h6F662074,
    32'h0A646E75,
    32'h00000000,
    32'h64616F4C,
    32'h20676E69,
    32'h6D6F7266,
    32'h49505320,
    32'h0000000A,
    32'h79706F43,
    32'h20676E69,
    32'h74736E49,
    32'h74637572,
    32'h736E6F69,
    32'h0000000A,
    32'h636F6C42,
    32'h0000206B,
    32'h6E6F6420,
    32'h00000A65,
    32'h79706F43,
    32'h20676E69,
    32'h61746144,
    32'h0000000A,
    32'h656E6F44,
    32'h756A202C,
    32'h6E69706D,
    32'h6F742067,
    32'h736E4920,
    32'h63757274,
    32'h6E6F6974,
    32'h4D415220,
    32'h00000A2E,
    32'h33323130,
    32'h37363534,
    32'h42413938,
    32'h46454443,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule