
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hEF410113,
    32'h00001D17,
    32'h9D0D0D13,
    32'h00001D97,
    32'h9C8D8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h00000513,
    32'h00000593,
    32'h014000EF,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'hCE86711D,
    32'h1080CCA2,
    32'h00EF4505,
    32'h45853C20,
    32'h00EF4501,
    32'h26236E20,
    32'hA039FE04,
    32'h27830001,
    32'h0785FEC4,
    32'hFEF42623,
    32'hFEC42703,
    32'h87936785,
    32'hD5E3BB77,
    32'h27B7FEE7,
    32'h07911A10,
    32'hC3984711,
    32'h262000EF,
    32'hCB8987AA,
    32'h02400593,
    32'h851367A5,
    32'h00EFA3C7,
    32'hA0017620,
    32'h67A545C5,
    32'hA6478513,
    32'h754000EF,
    32'h46014681,
    32'h451945A1,
    32'h414000EF,
    32'h00EF4501,
    32'h45814EE0,
    32'h00EF4505,
    32'h000154E0,
    32'h5A4000EF,
    32'h67C1872A,
    32'h8F7D17FD,
    32'h19E34785,
    32'h0693FEF7,
    32'h07B70200,
    32'h86138000,
    32'h45A13487,
    32'h07100513,
    32'h3DC000EF,
    32'h00EF4501,
    32'h45814B60,
    32'h00EF4505,
    32'h00015160,
    32'h56C000EF,
    32'h67C1872A,
    32'h8F7D17FD,
    32'h19E34785,
    32'h2423FEF7,
    32'h4581FE04,
    32'h00EF4521,
    32'h278343E0,
    32'h07A2FE84,
    32'h02000693,
    32'h45A1863E,
    32'h0EB00513,
    32'h398000EF,
    32'h10000513,
    32'h470000EF,
    32'h45094581,
    32'h4D0000EF,
    32'hFA040793,
    32'h10000593,
    32'h00EF853E,
    32'h278354A0,
    32'h2A23FA04,
    32'h2783FCF4,
    32'h2223FA44,
    32'h2783FEF4,
    32'h2823FA84,
    32'h2783FCF4,
    32'h2623FAC4,
    32'h2783FCF4,
    32'h2423FB04,
    32'h2783FCF4,
    32'h2023FB44,
    32'h2783FEF4,
    32'h2223FB84,
    32'h2783FCF4,
    32'h2023FBC4,
    32'h45D5FCF4,
    32'h851367A5,
    32'h00EFA787,
    32'h27836620,
    32'h2423FD44,
    32'h4581FEF4,
    32'h00EF4521,
    32'h2E233AE0,
    32'hA8B1FC04,
    32'hFE842783,
    32'h069307A2,
    32'h863E0200,
    32'h051345A1,
    32'h00EF0EB0,
    32'h65213020,
    32'h3DC000EF,
    32'h45094581,
    32'h43C000EF,
    32'h250365A1,
    32'h00EFFE44,
    32'h27034BA0,
    32'h6785FE44,
    32'h222397BA,
    32'h2703FEF4,
    32'h6785FE84,
    32'h242397BA,
    32'h2783FEF4,
    32'h853EFDC4,
    32'h1A6000EF,
    32'hFDC42783,
    32'h2E230785,
    32'h2703FCF4,
    32'h2783FDC4,
    32'h4FE3FCC4,
    32'h0001F8F7,
    32'h450000EF,
    32'h67C1872A,
    32'h8F7D17FD,
    32'h19E34785,
    32'h45B5FEF7,
    32'h851367A5,
    32'h00EFA907,
    32'h00EF5C60,
    32'h27836560,
    32'h2423FC84,
    32'h4581FEF4,
    32'h00EF4521,
    32'h2C2330E0,
    32'hA8B1FC04,
    32'hFE842783,
    32'h069307A2,
    32'h863E0200,
    32'h051345A1,
    32'h00EF0EB0,
    32'h65212620,
    32'h33C000EF,
    32'h45094581,
    32'h39C000EF,
    32'h250365A1,
    32'h00EFFE04,
    32'h270341A0,
    32'h6785FE04,
    32'h202397BA,
    32'h2703FEF4,
    32'h6785FE84,
    32'h242397BA,
    32'h2783FEF4,
    32'h853EFD84,
    32'h106000EF,
    32'hFD842783,
    32'h2C230785,
    32'h2703FCF4,
    32'h2783FD84,
    32'h4FE3FC04,
    32'h0593F8F7,
    32'h67A50220,
    32'hAA078513,
    32'h538000EF,
    32'h5C8000EF,
    32'h1A1077B7,
    32'hA02307A1,
    32'h05130007,
    32'h00EF0800,
    32'h47810AC0,
    32'h40F6853E,
    32'h61254466,
    32'h11018082,
    32'hCC22CE06,
    32'h26231000,
    32'h4681FE04,
    32'h45A14601,
    32'h09F00513,
    32'h1C8000EF,
    32'h04000513,
    32'h2A0000EF,
    32'h45014581,
    32'h248000EF,
    32'h45014581,
    32'h2F8000EF,
    32'hFE440793,
    32'h04000593,
    32'h00EF853E,
    32'h27833720,
    32'hD713FE44,
    32'h47850187,
    32'h00F70763,
    32'hFEC42783,
    32'h26230785,
    32'h2783FEF4,
    32'hD713FE44,
    32'h67C14087,
    32'h8F7D17FD,
    32'h21900793,
    32'h02F70263,
    32'hFE442783,
    32'h4087D713,
    32'h17FD67C1,
    32'h67898F7D,
    32'h076307E1,
    32'h278300F7,
    32'h0785FEC4,
    32'hFEF42623,
    32'hFEC42783,
    32'h40F2853E,
    32'h61054462,
    32'h11018082,
    32'h1000CE22,
    32'hFEA42623,
    32'hFEC42783,
    32'h00078067,
    32'h00010001,
    32'h00010001,
    32'h61054472,
    32'h71798082,
    32'hD422D606,
    32'h2E231800,
    32'h2783FCA4,
    32'h8BBDFDC4,
    32'hFEF42623,
    32'hFDC42783,
    32'h24238391,
    32'h4599FEF4,
    32'h851367A5,
    32'h00EFAC47,
    32'h270342E0,
    32'h67A5FE84,
    32'hAD478793,
    32'h458597BA,
    32'h00EF853E,
    32'h270341A0,
    32'h67A5FEC4,
    32'hAD478793,
    32'h458597BA,
    32'h00EF853E,
    32'h45994060,
    32'h851367A5,
    32'h00EFACC7,
    32'h00EF3FA0,
    32'h000148A0,
    32'h542250B2,
    32'h80826145,
    32'hFE010113,
    32'h00112E23,
    32'h00812C23,
    32'h02010413,
    32'hFEA42623,
    32'h00000593,
    32'h00F00513,
    32'h494000EF,
    32'h00000593,
    32'h00E00513,
    32'h488000EF,
    32'h00000593,
    32'h00D00513,
    32'h47C000EF,
    32'h00000593,
    32'h00C00513,
    32'h470000EF,
    32'hFEC42783,
    32'h00F05863,
    32'h00000593,
    32'h01000513,
    32'h45C000EF,
    32'hFEC42703,
    32'h00100793,
    32'h00E7D863,
    32'h00000593,
    32'h00B00513,
    32'h444000EF,
    32'hFEC42703,
    32'h00200793,
    32'h00E7D863,
    32'h00000593,
    32'h00000513,
    32'h42C000EF,
    32'hFEC42703,
    32'h00300793,
    32'h00E7D863,
    32'h00000593,
    32'h00100513,
    32'h414000EF,
    32'h00000013,
    32'h01C12083,
    32'h01812403,
    32'h02010113,
    32'h00008067,
    32'hFD010113,
    32'h02812623,
    32'h03010413,
    32'hFCA42E23,
    32'hFCB42C23,
    32'hFCC42A23,
    32'hFCD42823,
    32'h02000713,
    32'hFD842783,
    32'h40F707B3,
    32'hFDC42703,
    32'h00F717B3,
    32'hFEF42623,
    32'h1A1027B7,
    32'h00878793,
    32'hFEC42703,
    32'h00E7A023,
    32'h1A1027B7,
    32'h00C78793,
    32'hFD442703,
    32'h00E7A023,
    32'h1A1027B7,
    32'h01078793,
    32'hFD842703,
    32'h03F77693,
    32'hFD042703,
    32'h00871613,
    32'h00004737,
    32'hF0070713,
    32'h00E67733,
    32'h00E6E733,
    32'h00E7A023,
    32'h00000013,
    32'h02C12403,
    32'h03010113,
    32'h00008067,
    32'hFE010113,
    32'h00812E23,
    32'h02010413,
    32'hFEA42623,
    32'hFEB42423,
    32'h1A1027B7,
    32'h01478793,
    32'hFE842703,
    32'h01071713,
    32'h00070613,
    32'hFEC42683,
    32'h00010737,
    32'hFFF70713,
    32'h00E6F733,
    32'h00E66733,
    32'h00E7A023,
    32'h00000013,
    32'h01C12403,
    32'h02010113,
    32'h00008067,
    32'hFD010113,
    32'h02812623,
    32'h03010413,
    32'hFCA42E23,
    32'h1A1027B7,
    32'h01078793,
    32'h0007A783,
    32'hFEF42623,
    32'hFDC42783,
    32'h01079793,
    32'h00078713,
    32'hFEC42783,
    32'h00078693,
    32'h000107B7,
    32'hFFF78793,
    32'h00F6F7B3,
    32'h00F767B3,
    32'hFEF42623,
    32'h1A1027B7,
    32'h01078793,
    32'hFEC42703,
    32'h00E7A023,
    32'h00000013,
    32'h02C12403,
    32'h03010113,
    32'h00008067,
    32'hFE010113,
    32'h00812E23,
    32'h02010413,
    32'hFEA42623,
    32'hFEB42423,
    32'h1A1027B7,
    32'hFE842703,
    32'h00870713,
    32'h00100693,
    32'h00E696B3,
    32'h00001737,
    32'hF0070713,
    32'h00E6F6B3,
    32'h00100613,
    32'hFEC42703,
    32'h00E61733,
    32'h0FF77713,
    32'h00E6E733,
    32'h00E7A023,
    32'h00000013,
    32'h01C12403,
    32'h02010113,
    32'h00008067,
    32'hFE010113,
    32'h00812E23,
    32'h02010413,
    32'h1A1027B7,
    32'h0007A783,
    32'hFEF42623,
    32'hFEC42783,
    32'h00078513,
    32'h01C12403,
    32'h02010113,
    32'h00008067,
    32'hFD010113,
    32'h02812623,
    32'h03010413,
    32'hFCA42E23,
    32'hFCB42C23,
    32'hFD842783,
    32'h4057D793,
    32'h7FF7F793,
    32'hFEF42623,
    32'hFD842783,
    32'h01F7F793,
    32'h00078863,
    32'hFEC42783,
    32'h00178793,
    32'hFEF42623,
    32'hFE042423,
    32'h0480006F,
    32'h00000013,
    32'h1A1027B7,
    32'h0007A783,
    32'h4107D793,
    32'h0FF7F793,
    32'hFE0788E3,
    32'hFE842783,
    32'h00279793,
    32'hFDC42703,
    32'h00F707B3,
    32'h1A102737,
    32'h02070713,
    32'h00072703,
    32'h00E7A023,
    32'hFE842783,
    32'h00178793,
    32'hFEF42423,
    32'hFE842703,
    32'hFEC42783,
    32'hFAF74AE3,
    32'h00000013,
    32'h02C12403,
    32'h03010113,
    32'h00008067,
    32'hFE010113,
    32'h00812E23,
    32'h02010413,
    32'hFEA42623,
    32'h00058793,
    32'hFEF41523,
    32'h1A1077B7,
    32'h00478793,
    32'h1A107737,
    32'h00470713,
    32'h00072703,
    32'h00276713,
    32'h00E7A023,
    32'h1A1007B7,
    32'h00C78793,
    32'h08300713,
    32'h00E7A023,
    32'h1A1007B7,
    32'h00478793};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule