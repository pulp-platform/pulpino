
`define RISCV
