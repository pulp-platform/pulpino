
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h81868106,
    32'h82868206,
    32'h83868306,
    32'h84868406,
    32'h85868506,
    32'h86868606,
    32'h87868706,
    32'h88868806,
    32'h89868906,
    32'h8A868A06,
    32'h8B868B06,
    32'h8C868C06,
    32'h8D868D06,
    32'h8E868E06,
    32'h8F868F06,
    32'h00100117,
    32'hF3010113,
    32'h00000D17,
    32'h5D8D0D13,
    32'h00000D97,
    32'h5D0D8D93,
    32'h01BD5763,
    32'h000D2023,
    32'hDDE30D11,
    32'h0513FFAD,
    32'h05930000,
    32'h00EF0000,
    32'h00000740,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h11010000,
    32'h46014681,
    32'h051345A1,
    32'hCE0609F0,
    32'h348000EF,
    32'h04000513,
    32'h384000EF,
    32'h45014581,
    32'h36C000EF,
    32'h45014581,
    32'h394000EF,
    32'h05930028,
    32'h00EF0400,
    32'h47A23BE0,
    32'h21900713,
    32'h0187D513,
    32'h157D87A1,
    32'h1007D7B3,
    32'h00A03533,
    32'h00E78863,
    32'h07616709,
    32'h37B38F99,
    32'h953E00F0,
    32'h610540F2,
    32'h715D8082,
    32'hC6864505,
    32'hC2A6C4A2,
    32'hDE4EC0CA,
    32'hDA56DC52,
    32'hD65ED85A,
    32'hD266D462,
    32'h00EFD06A,
    32'h45852660,
    32'h00EF4501,
    32'h67853BA0,
    32'hBB878793,
    32'h0037C0FB,
    32'h00010001,
    32'h27B74711,
    32'hC3D81A10,
    32'hF63FF0EF,
    32'h8537C911,
    32'h05930000,
    32'h05130240,
    32'h00EF6085,
    32'hA0013DA0,
    32'h00008537,
    32'h051345C5,
    32'h00EF6305,
    32'h46813CA0,
    32'h45A14601,
    32'h00EF4519,
    32'h450128A0,
    32'h2C8000EF,
    32'h458164C1,
    32'h00EF4505,
    32'h14FD2DE0,
    32'h00EF4405,
    32'h8D652FA0,
    32'hFE851DE3,
    32'h80000637,
    32'h02000693,
    32'h34860613,
    32'h051345A1,
    32'h00EF0710,
    32'h45012560,
    32'h294000EF,
    32'h458164C1,
    32'h00EF8522,
    32'h14FD2AA0,
    32'h2C8000EF,
    32'h1DE38D65,
    32'h4581FE85,
    32'h00EF4521,
    32'h06932660,
    32'h46010200,
    32'h051345A1,
    32'h00EF0EB0,
    32'h05132220,
    32'h00EF1000,
    32'h458125E0,
    32'h00EF4509,
    32'h05932760,
    32'h850A1000,
    32'h2A0000EF,
    32'h00008537,
    32'h45D54CB2,
    32'h64450513,
    32'h4C124402,
    32'h4AD249C2,
    32'h00EF4B72,
    32'h45813220,
    32'h00EF4521,
    32'h5F6321A0,
    32'h84A20790,
    32'h49016421,
    32'h409C0C33,
    32'h00008BB7,
    32'h6A040413,
    32'h00008A37,
    32'h96136D05,
    32'h06930084,
    32'h45A10200,
    32'h0EB00513,
    32'h1B8000EF,
    32'h00EF6521,
    32'h45811F60,
    32'h00EF4509,
    32'h053320E0,
    32'h65A1009C,
    32'h238000EF,
    32'h85134599,
    32'h00EF65CB,
    32'h55132CA0,
    32'h45850049,
    32'h00EF9522,
    32'h75132BE0,
    32'h458500F9,
    32'h00EF9522,
    32'h09052B20,
    32'h05134599,
    32'h00EF664A,
    32'h94EA2A60,
    32'h2CC000EF,
    32'hFB2C91E3,
    32'h147D6441,
    32'h00EF4485,
    32'h8D611E60,
    32'hFE951DE3,
    32'h00008537,
    32'h051345B5,
    32'h00EF66C5,
    32'h00EF27E0,
    32'h45812A60,
    32'h00EF4521,
    32'h5F631720,
    32'h64210760,
    32'h490184CE,
    32'h413A89B3,
    32'h00008BB7,
    32'h6A040413,
    32'h00008A37,
    32'h96136A85,
    32'h06930084,
    32'h45A10200,
    32'h0EB00513,
    32'h110000EF,
    32'h00EF6521,
    32'h458114E0,
    32'h00EF4509,
    32'h85331660,
    32'h65A10099,
    32'h190000EF,
    32'h85134599,
    32'h00EF65CB,
    32'h55132220,
    32'h45850049,
    32'h00EF9522,
    32'h75132160,
    32'h458500F9,
    32'h00EF9522,
    32'h090520A0,
    32'h05134599,
    32'h00EF664A,
    32'h94D61FE0,
    32'h224000EF,
    32'hFB2B11E3,
    32'h00008537,
    32'h02200593,
    32'h67C50513,
    32'h1E4000EF,
    32'h20C000EF,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000793,
    32'h00078067,
    32'h00010001,
    32'h40B60001,
    32'h44264501,
    32'h49064496,
    32'h5A6259F2,
    32'h5B425AD2,
    32'h5C225BB2,
    32'h5D025C92,
    32'h80826161,
    32'hC4221141,
    32'h842A4581,
    32'hC606453D,
    32'h00EFC226,
    32'h45811D60,
    32'h00EF4539,
    32'h45811CE0,
    32'h00EF4535,
    32'h45811C60,
    32'h00EF4531,
    32'h5F631BE0,
    32'h44850280,
    32'h45414581,
    32'h1B0000EF,
    32'h02940863,
    32'h452D4581,
    32'h1A4000EF,
    32'h01634789,
    32'h458102F4,
    32'h00EF4501,
    32'h478D1960,
    32'h00F40A63,
    32'h40B28526,
    32'h44924422,
    32'h01414581,
    32'h1800006F,
    32'h442240B2,
    32'h01414492,
    32'h00008082,
    32'h08136811,
    32'h06A2F008,
    32'h02000713,
    32'h1A1027B7,
    32'hF6B38F0D,
    32'hF5930106,
    32'h153303F5,
    32'h881300E5,
    32'h87130087,
    32'h8DD500C7,
    32'h202307C1,
    32'hC31000A8,
    32'h8082C38C,
    32'h553305C2,
    32'h8DC91005,
    32'h1A1027B7,
    32'h8082CBCC,
    32'h1A102737,
    32'h431C0741,
    32'hC63E1141,
    32'h054247B2,
    32'h1007D7B3,
    32'hC62A8D5D,
    32'h014147B2,
    32'h8082C31C,
    32'h05A14785,
    32'h00B795B3,
    32'h00A79533,
    32'h87936785,
    32'h8DFDF007,
    32'h0FF57513,
    32'h27B78D4D,
    32'hC3881A10,
    32'h00008082,
    32'h1A1027B7,
    32'h1141439C,
    32'h4532C63E,
    32'h80820141,
    32'h4055D793,
    32'hF7931141,
    32'h89FD7FF7,
    32'hC581C43E,
    32'h078547A2,
    32'hC602C43E,
    32'h47A246B2,
    32'h1A102737,
    32'h02070813,
    32'h02F6D463,
    32'h87C1431C,
    32'h0FF7F793,
    32'h47B2DFE5,
    32'h00082583,
    32'h078A46B2,
    32'hC6360685,
    32'h46A24632,
    32'h1EB56023,
    32'hFED640E3,
    32'h80820141,
    32'h1A107737,
    32'h43100711,
    32'h1A1007B7,
    32'h00266613,
    32'h8513C310,
    32'h071300C7,
    32'hC1180830,
    32'h00478693,
    32'h0085D813,
    32'hF5934721,
    32'hA0230FF5,
    32'hE02B0106,
    32'h07131CB7,
    32'hC3980A70,
    32'hC11C478D,
    32'hF793429C,
    32'hE7930F07,
    32'hC29C0027,
    32'h00008082,
    32'h1A100737,
    32'hC1850751,
    32'h04000693,
    32'hF793431C,
    32'hDFED0207,
    32'h0015460B,
    32'h1A1007B7,
    32'hC39015FD,
    32'hE29916FD,
    32'h8082F1F5,
    32'h8082F1F5,
    32'h1A100737,
    32'h431C0751,
    32'h0407F793,
    32'h8082DFED,
    32'h1A1076B7,
    32'h1141429C,
    32'h4785C63E,
    32'h97B34732,
    32'hC79300A7,
    32'h8FF9FFF7,
    32'h47B2C63E,
    32'h00A595B3,
    32'h00F5E533,
    32'h47B2C62A,
    32'hC29C0141,
    32'h00008082,
    32'h4F525245,
    32'h53203A52,
    32'h736E6170,
    32'h206E6F69,
    32'h20495053,
    32'h73616C66,
    32'h6F6E2068,
    32'h6F662074,
    32'h0A646E75,
    32'h00000000,
    32'h64616F4C,
    32'h20676E69,
    32'h6D6F7266,
    32'h49505320,
    32'h0000000A,
    32'h79706F43,
    32'h20676E69,
    32'h74736E49,
    32'h74637572,
    32'h736E6F69,
    32'h0000000A,
    32'h636F6C42,
    32'h0000206B,
    32'h6E6F6420,
    32'h00000A65,
    32'h79706F43,
    32'h20676E69,
    32'h61746144,
    32'h0000000A,
    32'h656E6F44,
    32'h756A202C,
    32'h6E69706D,
    32'h6F742067,
    32'h736E4920,
    32'h63757274,
    32'h6E6F6974,
    32'h4D415220,
    32'h00000A2E,
    32'h33323130,
    32'h37363534,
    32'h42413938,
    32'h46454443,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule