`define PULP_FPGA_EMUL

//`define RISCV
