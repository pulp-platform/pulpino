//`define SHARED_APU
`define APU