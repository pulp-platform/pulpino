
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:699] [31:0] mem = {
    32'h0040006F,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hF8010113,
    32'h00001D17,
    32'h918D0D13,
    32'h00001D97,
    32'h910D8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h00000513,
    32'h00000593,
    32'h0A0000EF,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'hFE010113,
    32'h00000693,
    32'h00000613,
    32'h00800593,
    32'h09F00513,
    32'h00112E23,
    32'h48C000EF,
    32'h04000513,
    32'h4D8000EF,
    32'h00000593,
    32'h00000513,
    32'h4B0000EF,
    32'h00000593,
    32'h00000513,
    32'h4F8000EF,
    32'h00810513,
    32'h04000593,
    32'h538000EF,
    32'h00812783,
    32'h21900713,
    32'h0187D513,
    32'h4087D793,
    32'h01079793,
    32'hFFF50513,
    32'h0107D793,
    32'h00A03533,
    32'h00E78C63,
    32'h00002737,
    32'h01870713,
    32'h40E787B3,
    32'h00F037B3,
    32'h00F50533,
    32'h01C12083,
    32'h02010113,
    32'h00008067,
    32'hFB010113,
    32'h00100513,
    32'h04112623,
    32'h04812423,
    32'h04912223,
    32'h05212023,
    32'h03312E23,
    32'h03412C23,
    32'h03512A23,
    32'h03612823,
    32'h03712623,
    32'h03812423,
    32'h03912223,
    32'h03A12023,
    32'h32C000EF,
    32'h00100593,
    32'h00000513,
    32'h52C000EF,
    32'h000017B7,
    32'hBB878793,
    32'h00000013,
    32'hFFF78793,
    32'hFE079CE3,
    32'h00400713,
    32'h1A1027B7,
    32'h00E7A223,
    32'hF0DFF0EF,
    32'h00050C63,
    32'h00008537,
    32'h02400593,
    32'h7A850513,
    32'h544000EF,
    32'h0000006F,
    32'h00008537,
    32'h01100593,
    32'h7D050513,
    32'h530000EF,
    32'h00000693,
    32'h00000613,
    32'h00800593,
    32'h00600513,
    32'h374000EF,
    32'h00000513,
    32'h3C0000EF,
    32'h000104B7,
    32'h00000593,
    32'h00100513,
    32'h3E8000EF,
    32'hFFF48493,
    32'h00100413,
    32'h40C000EF,
    32'h00957533,
    32'hFE851CE3,
    32'h80000637,
    32'h02000693,
    32'h34860613,
    32'h00800593,
    32'h07100513,
    32'h330000EF,
    32'h00000513,
    32'h37C000EF,
    32'h000104B7,
    32'h00000593,
    32'h00040513,
    32'h3A4000EF,
    32'hFFF48493,
    32'h3CC000EF,
    32'h00957533,
    32'hFE851CE3,
    32'h00000593,
    32'h00800513,
    32'h334000EF,
    32'h02000693,
    32'h00000613,
    32'h00800593,
    32'h0EB00513,
    32'h2E8000EF,
    32'h10000513,
    32'h334000EF,
    32'h00000593,
    32'h00200513,
    32'h360000EF,
    32'h10000593,
    32'h00010513,
    32'h3A0000EF,
    32'h00C12C83,
    32'h00008537,
    32'h01500593,
    32'h7E450513,
    32'h00012403,
    32'h00412C03,
    32'h01012983,
    32'h01412A83,
    32'h01C12B03,
    32'h448000EF,
    32'h00000593,
    32'h00800513,
    32'h2CC000EF,
    32'h0B905063,
    32'h00040493,
    32'h00009437,
    32'h00000913,
    32'h409C0C33,
    32'h00008BB7,
    32'h84040413,
    32'h00009A37,
    32'h00001D37,
    32'h00849613,
    32'h02000693,
    32'h00800593,
    32'h0EB00513,
    32'h25C000EF,
    32'h00008537,
    32'h2A8000EF,
    32'h00000593,
    32'h00200513,
    32'h2D4000EF,
    32'h009C0533,
    32'h000085B7,
    32'h314000EF,
    32'h00600593,
    32'h7FCB8513,
    32'h3D8000EF,
    32'h00495513,
    32'h00100593,
    32'h00A40533,
    32'h3C8000EF,
    32'h00F97513,
    32'h00100593,
    32'h00A40533,
    32'h3B8000EF,
    32'h00190913,
    32'h00600593,
    32'h804A0513,
    32'h3A8000EF,
    32'h01A484B3,
    32'h3DC000EF,
    32'hF92C94E3,
    32'h00010437,
    32'hFFF40413,
    32'h00100493,
    32'h2A0000EF,
    32'h00857533,
    32'hFE951CE3,
    32'h00009537,
    32'h00D00593,
    32'h80C50513,
    32'h374000EF,
    32'h3AC000EF,
    32'h00000593,
    32'h00800513,
    32'h1F4000EF,
    32'h0B605063,
    32'h00009437,
    32'h00098493,
    32'h00000913,
    32'h413A89B3,
    32'h00008BB7,
    32'h84040413,
    32'h00009A37,
    32'h00001AB7,
    32'h00849613,
    32'h02000693,
    32'h00800593,
    32'h0EB00513,
    32'h184000EF,
    32'h00008537,
    32'h1D0000EF,
    32'h00000593,
    32'h00200513,
    32'h1FC000EF,
    32'h00998533,
    32'h000085B7,
    32'h23C000EF,
    32'h00600593,
    32'h7FCB8513,
    32'h300000EF,
    32'h00495513,
    32'h00100593,
    32'h00A40533,
    32'h2F0000EF,
    32'h00F97513,
    32'h00100593,
    32'h00A40533,
    32'h2E0000EF,
    32'h00190913,
    32'h00600593,
    32'h804A0513,
    32'h2D0000EF,
    32'h015484B3,
    32'h304000EF,
    32'hF92B14E3,
    32'h00009537,
    32'h02200593,
    32'h81C50513,
    32'h2B4000EF,
    32'h2EC000EF,
    32'h08000793,
    32'h00078067,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h04C12083,
    32'h00000513,
    32'h04812403,
    32'h04412483,
    32'h04012903,
    32'h03C12983,
    32'h03812A03,
    32'h03412A83,
    32'h03012B03,
    32'h02C12B83,
    32'h02812C03,
    32'h02412C83,
    32'h02012D03,
    32'h05010113,
    32'h00008067,
    32'hFF010113,
    32'h00812423,
    32'h00000593,
    32'h00050413,
    32'h00F00513,
    32'h00112623,
    32'h00912223,
    32'h290000EF,
    32'h00000593,
    32'h00E00513,
    32'h284000EF,
    32'h00000593,
    32'h00D00513,
    32'h278000EF,
    32'h00000593,
    32'h00C00513,
    32'h26C000EF,
    32'h04805E63,
    32'h00100493,
    32'h00000593,
    32'h01000513,
    32'h258000EF,
    32'h04940463,
    32'h00000593,
    32'h00B00513,
    32'h248000EF,
    32'h00200793,
    32'h02F40A63,
    32'h00000593,
    32'h00000513,
    32'h234000EF,
    32'h00300793,
    32'h02F40063,
    32'h00048513,
    32'h00C12083,
    32'h00812403,
    32'h00412483,
    32'h00000593,
    32'h01010113,
    32'h2100006F,
    32'h00C12083,
    32'h00812403,
    32'h00412483,
    32'h01010113,
    32'h00008067,
    32'h00004737,
    32'hF0070713,
    32'h00869693,
    32'h02000793,
    32'h40B787B3,
    32'h00E6F6B3,
    32'h03F5F593,
    32'h1A102737,
    32'h00F51533,
    32'h00B6E5B3,
    32'h00A72423,
    32'h00C72623,
    32'h00B72823,
    32'h00008067,
    32'h01051513,
    32'h01059593,
    32'h01055513,
    32'h00A5E5B3,
    32'h1A1027B7,
    32'h00B7AA23,
    32'h00008067,
    32'h1A102737,
    32'h01072783,
    32'hFF010113,
    32'h01051513,
    32'h00F12623,
    32'h00C12783,
    32'h01079793,
    32'h0107D793,
    32'h00F56533,
    32'h00A12623,
    32'h00C12783,
    32'h01010113,
    32'h00F72823,
    32'h00008067,
    32'h00100793,
    32'h00858593,
    32'h00B795B3,
    32'h00A79533,
    32'h000017B7,
    32'hF0078793,
    32'h00F5F5B3,
    32'h0FF57513,
    32'h00A5E533,
    32'h1A1027B7,
    32'h00A7A023,
    32'h00008067,
    32'h1A1027B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12503,
    32'h01010113,
    32'h00008067,
    32'h4055D793,
    32'hFF010113,
    32'h7FF7F793,
    32'h01F5F593,
    32'h00F12423,
    32'h00058863,
    32'h00812783,
    32'h00178793,
    32'h00F12423,
    32'h00012623,
    32'h00C12683,
    32'h00812783,
    32'h1A102737,
    32'h00070813,
    32'h04F6D063,
    32'h00072783,
    32'h4107D793,
    32'h0FF7F793,
    32'hFE078AE3,
    32'h00C12783,
    32'h02082583,
    32'h00C12683,
    32'h00279793,
    32'h00F507B3,
    32'h00168693,
    32'h00D12623,
    32'h00C12603,
    32'h00812683,
    32'h00B7A023,
    32'hFCD644E3,
    32'h01010113,
    32'h00008067,
    32'h1A1076B7,
    32'h0046A703,
    32'h1A1007B7,
    32'h0085D613,
    32'h00276713,
    32'h00E6A223,
    32'h08300713,
    32'h00E7A623,
    32'h0FF5F593,
    32'h0A700713,
    32'h00C7A223,
    32'h00B7A023,
    32'h00E7A423,
    32'h00300713,
    32'h00E7A623,
    32'h0047A703,
    32'h0F077713,
    32'h00276713,
    32'h00E7A223,
    32'h00008067,
    32'h1A100737,
    32'h02058A63,
    32'h04050613,
    32'h01472783,
    32'h0207F793,
    32'hFE078CE3,
    32'h00150513,
    32'hFFF54683,
    32'h1A1007B7,
    32'hFFF58593,
    32'h00D7A023,
    32'hFCC50CE3,
    32'hFC059EE3,
    32'h00008067,
    32'h00008067,
    32'h1A100737,
    32'h01472783,
    32'h0407F793,
    32'hFE078CE3,
    32'h00008067,
    32'h1A1076B7,
    32'h0006A783,
    32'hFF010113,
    32'h00A595B3,
    32'h00F12623,
    32'h00C12703,
    32'h00100793,
    32'h00A797B3,
    32'hFFF7C793,
    32'h00E7F7B3,
    32'h00F12623,
    32'h00C12783,
    32'h00F5E533,
    32'h00A12623,
    32'h00C12783,
    32'h01010113,
    32'h00F6A023,
    32'h00008067,
    32'h4F525245,
    32'h53203A52,
    32'h736E6170,
    32'h206E6F69,
    32'h20495053,
    32'h73616C66,
    32'h6F6E2068,
    32'h6F662074,
    32'h0A646E75,
    32'h00000000,
    32'h64616F4C,
    32'h20676E69,
    32'h6D6F7266,
    32'h49505320,
    32'h0000000A,
    32'h79706F43,
    32'h20676E69,
    32'h74736E49,
    32'h74637572,
    32'h736E6F69,
    32'h0000000A,
    32'h636F6C42,
    32'h0000206B,
    32'h6E6F6420,
    32'h00000A65,
    32'h79706F43,
    32'h20676E69,
    32'h61746144,
    32'h0000000A,
    32'h656E6F44,
    32'h756A202C,
    32'h6E69706D,
    32'h6F742067,
    32'h736E4920,
    32'h63757274,
    32'h6E6F6974,
    32'h4D415220,
    32'h00000A2E,
    32'h33323130,
    32'h37363534,
    32'h42413938,
    32'h46454443,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000014,
    32'h00000018,
    32'hFFFFF858,
    32'h0000008C,
    32'h200E4400,
    32'h7F011154,
    32'h00000038,
    32'h00000030,
    32'hFFFFF8CC,
    32'h00000364,
    32'h500E4400,
    32'h7F011174,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h117A1411,
    32'h16117915,
    32'h77171178,
    32'h11761811,
    32'h1A117519,
    32'h00000074,
    32'h0000001C,
    32'h0000006C,
    32'hFFFFFBF4,
    32'h000000B4,
    32'h100E4400,
    32'h7E081148,
    32'h7F011150,
    32'h007D0911,
    32'h00000010,
    32'h0000008C,
    32'hFFFFFC88,
    32'h00000038,
    32'h00000000,
    32'h00000010,
    32'h000000A0,
    32'hFFFFFCAC,
    32'h0000001C,
    32'h00000000,
    32'h00000010,
    32'h000000B4,
    32'hFFFFFCB4,
    32'h00000038,
    32'h100E4C00,
    32'h00000010,
    32'h000000C8,
    32'hFFFFFCD8,
    32'h00000030,
    32'h00000000,
    32'h00000010,
    32'h000000DC,
    32'hFFFFFCF4,
    32'h0000001C,
    32'h100E4C00,
    32'h00000010,
    32'h000000F0,
    32'hFFFFFCFC,
    32'h00000080,
    32'h100E4800,
    32'h00000010,
    32'h00000104,
    32'hFFFFFD68,
    32'h00000050,
    32'h00000000,
    32'h00000010,
    32'h00000118,
    32'hFFFFFDA4,
    32'h0000003C,
    32'h00000000,
    32'h00000010,
    32'h0000012C,
    32'hFFFFFDCC,
    32'h00000014,
    32'h00000000,
    32'h00000010,
    32'h00000140,
    32'hFFFFFDCC,
    32'h00000048,
    32'h100E4C00,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule